entity scalar is
end entity;

architecture test of scalar is
    signal x : integer;
begin

    process is
    begin
        x <= 1;
    end process;

end architecture;
